	double geophysical_variable(time) ;
		geophysical_variable:_FillValue = -999. ;
		geophysical_variable:accuracy = " " ;
		geophysical_variable:ancillary_variables = "geophysical_variable_qc" ;
		geophysical_variable:instrument = " " ;
		geophysical_variable:long_name = " " ;
		geophysical_variable:observation_type = " " ;
		geophysical_variable:platform = "platform" ;
		geophysical_variable:precision = " " ;
		geophysical_variable:resolution = " " ;
		geophysical_variable:standard_name = " " ;
		geophysical_variable:units = " " ;
		geophysical_variable:valid_max = 40. ;
		geophysical_variable:valid_min = -5. ;
	byte geophysical_variable_qc(time) ;
		geophysical_variable_qc:_FillValue = -127b ;
		geophysical_variable_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed not_used not_used interpolated_value missing_value" ;
		geophysical_variable_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		geophysical_variable_qc:long_name = "geophysical_variable Quality Flag" ;
		geophysical_variable_qc:standard_name = "geophysical_variable status_flag" ;
		geophysical_variable_qc:valid_max = 9b ;
		geophysical_variable_qc:valid_min = 0b ;
