netcdf IOOS_Glider_NetCDF_v3.0-noqartod {
dimensions:
	time = UNLIMITED ; // (0 currently)
	traj_strlen = 20 ;
variables:
	double conductivity(time) ;
		conductivity:_FillValue = -999. ;
		conductivity:accuracy = " " ;
		conductivity:ancillary_variables = " " ;
		conductivity:instrument = "instrument_ctd" ;
		conductivity:long_name = "Conductivity" ;
		conductivity:observation_type = "measured" ;
		conductivity:platform = "platform" ;
		conductivity:precision = " " ;
		conductivity:resolution = " " ;
		conductivity:standard_name = "sea_water_electrical_conductivity" ;
		conductivity:units = "S m-1" ;
		conductivity:valid_max = 10. ;
		conductivity:valid_min = 0. ;
	double density(time) ;
		density:_FillValue = -999. ;
		density:accuracy = " " ;
		density:ancillary_variables = " " ;
		density:instrument = "instrument_ctd" ;
		density:long_name = "Density" ;
		density:observation_type = "calculated" ;
		density:platform = "platform" ;
		density:precision = " " ;
		density:resolution = " " ;
		density:standard_name = "sea_water_density" ;
		density:units = "kg m-3" ;
		density:valid_max = 1040. ;
		density:valid_min = 1015. ;
	double depth(time) ;
		depth:_FillValue = -999. ;
		depth:accuracy = " " ;
		depth:ancillary_variables = " " ;
		depth:comment = " " ;
		depth:instrument = "instrument_ctd" ;
		depth:long_name = "Depth" ;
		depth:observation_type = "calculated" ;
		depth:platform = "platform" ;
		depth:positive = "down" ;
		depth:precision = " " ;
		depth:reference_datum = "sea-surface" ;
		depth:resolution = " " ;
		depth:standard_name = "depth" ;
		depth:units = "m" ;
		depth:valid_max = 2000 ;
		depth:valid_min = 0 ;
	int instrument_ctd ;
		instrument_ctd:_FillValue = -999 ;
		instrument_ctd:calibration_date = " " ;
		instrument_ctd:calibration_report = " " ;
		instrument_ctd:comment = "pumped CTD" ;
		instrument_ctd:factory_calibrated = " " ;
		instrument_ctd:long_name = "Seabird Glider Payload CTD" ;
		instrument_ctd:make_model = "Seabird GPCTD" ;
		instrument_ctd:platform = "platform" ;
		instrument_ctd:serial_number = " " ;
		instrument_ctd:type = "platform" ;
	double lat(time) ;
		lat:_FillValue = -999. ;
		lat:ancillary_variables = " " ;
		lat:comment = "Interpolated latitude at each point in the time-series" ;
		lat:coordinate_reference_frame = "urn:ogc:crs:EPSG::4326" ;
		lat:long_name = "Latitude" ;
		lat:observation_type = "measured" ;
		lat:platform = "platform" ;
		lat:reference = "WGS84" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:valid_max = 90. ;
		lat:valid_min = -90. ;
	double lat_uv ;
		lat_uv:_FillValue = -999. ;
		lat_uv:comment = "The depth-averaged current is an estimate of the net current measured while the glider is underwater.  The value is calculated over the entire underwater segment, which may consist of 1 or more dives." ;
		lat_uv:long_name = "Depth-Averaged Latitude" ;
		lat_uv:observation_type = "calculated" ;
		lat_uv:platform = "platform" ;
		lat_uv:standard_name = "latitude" ;
		lat_uv:units = "degrees_north" ;
		lat_uv:valid_max = 90. ;
		lat_uv:valid_min = -90. ;
	double lon(time) ;
		lon:_FillValue = -999. ;
		lon:ancillary_variables = " " ;
		lon:comment = "Interpolated longitude at each point in the time-series." ;
		lon:coordinate_reference_frame = "urn:ogc:crs:EPSG::4326" ;
		lon:long_name = "Longitude" ;
		lon:observation_type = "measured" ;
		lon:platform = "platform" ;
		lon:reference = "WGS84" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:valid_max = 180. ;
		lon:valid_min = -180. ;
	double lon_uv ;
		lon_uv:_FillValue = -999. ;
		lon_uv:comment = "The depth-averaged current is an estimate of the net current measured while the glider is underwater.  The value is calculated over the entire underwater segment, which may consist of 1 or more dives." ;
		lon_uv:long_name = "Depth-Averaged Longitude" ;
		lon_uv:observation_type = "calculated" ;
		lon_uv:platform = "platform" ;
		lon_uv:standard_name = "longitude" ;
		lon_uv:units = "degrees_east" ;
		lon_uv:valid_max = 180. ;
		lon_uv:valid_min = -180. ;
	int platform ;
		platform:_FillValue = -999 ;
		platform:comment = " " ;
		platform:id = " " ;
		platform:instrument = "instrument_ctd" ;
		platform:long_name = " " ;
		platform:type = "platform" ;
		platform:wmo_id = " " ;
	double pressure(time) ;
		pressure:_FillValue = -999. ;
		pressure:accuracy = " " ;
		pressure:ancillary_variables = " " ;
		pressure:comment = " " ;
		pressure:instrument = "instrument_ctd" ;
		pressure:long_name = "Pressure" ;
		pressure:observation_type = "measured" ;
		pressure:platform = "platform" ;
		pressure:positive = "down" ;
		pressure:precision = " " ;
		pressure:reference_datum = "sea-surface" ;
		pressure:resolution = " " ;
		pressure:standard_name = "sea_water_pressure" ;
		pressure:units = "dbar" ;
		pressure:valid_max = 2000 ;
		pressure:valid_min = 0 ;
	int profile_id ;
		profile_id:_FillValue = -999 ;
		profile_id:comment = "Sequential profile number within the trajectory.  This value is unique in each file that is part of a single trajectory/deployment." ;
		profile_id:long_name = "Profile ID" ;
		profile_id:valid_max = 2147483647 ;
		profile_id:valid_min = 1 ;
	double profile_lat ;
		profile_lat:_FillValue = -999. ;
		profile_lat:comment = "Value is interpolated to provide an estimate of the latitude at the mid-point of the profile" ;
		profile_lat:long_name = "Profile Center Latitude" ;
		profile_lat:observation_type = "calculated" ;
		profile_lat:platform = "platform" ;
		profile_lat:standard_name = "latitude" ;
		profile_lat:units = "degrees_north" ;
		profile_lat:valid_max = 90. ;
		profile_lat:valid_min = -90. ;
	double profile_lon ;
		profile_lon:_FillValue = -999. ;
		profile_lon:comment = "Value is interpolated to provide an estimate of the longitude at the mid-point of the profile" ;
		profile_lon:long_name = "Profile Center Longitude" ;
		profile_lon:observation_type = "calculated" ;
		profile_lon:platform = "platform" ;
		profile_lon:standard_name = "longitude" ;
		profile_lon:units = "degrees_east" ;
		profile_lon:valid_max = 180. ;
		profile_lon:valid_min = -180. ;
	double profile_time ;
		profile_time:_FillValue = -999. ;
		profile_time:calendar = "gregorian" ;
		profile_time:comment = "Timestamp corresponding to the mid-point of the profile" ;
		profile_time:long_name = "Profile Center Time" ;
		profile_time:observation_type = "calculated" ;
		profile_time:platform = "platform" ;
		profile_time:standard_name = "time" ;
		profile_time:units = "seconds since 1970-01-01T00:00:00Z" ;
	double salinity(time) ;
		salinity:_FillValue = -999. ;
		salinity:accuracy = " " ;
		salinity:ancillary_variables = " " ;
		salinity:instrument = "instrument_ctd" ;
		salinity:long_name = "Salinity" ;
		salinity:observation_type = "calculated" ;
		salinity:platform = "platform" ;
		salinity:precision = " " ;
		salinity:resolution = " " ;
		salinity:standard_name = "sea_water_practical_salinity" ;
		salinity:units = 1 ;
		salinity:valid_max = 40. ;
		salinity:valid_min = 0. ;
	double temperature(time) ;
		temperature:_FillValue = -999. ;
		temperature:accuracy = " " ;
		temperature:ancillary_variables = " " ;
		temperature:instrument = "instrument_ctd" ;
		temperature:long_name = "Temperature" ;
		temperature:observation_type = "measured" ;
		temperature:platform = "platform" ;
		temperature:precision = " " ;
		temperature:resolution = " " ;
		temperature:standard_name = "sea_water_temperature" ;
		temperature:units = "Celsius" ;
		temperature:valid_max = 40. ;
		temperature:valid_min = -5. ;
	double time(time) ;
		time:ancillary_variables = " " ;
		time:calendar = "gregorian" ;
		time:comment = "Measured or calculated time at each point in the time-series" ;
		time:long_name = "Time" ;
		time:observation_type = "measured" ;
		time:standard_name = "time" ;
		time:units = "seconds since 1970-01-01T00:00:00Z" ;
	double time_uv ;
		time_uv:_FillValue = -999. ;
		time_uv:calendar = "gregorian" ;
		time_uv:comment = "The depth-averaged current is an estimate of the net current measured while the glider is underwater.  The value is calculated over the entire underwater segment, which may consist of 1 or more dives." ;
		time_uv:long_name = "Depth-Averaged Time" ;
		time_uv:observation_type = "calculated" ;
		time_uv:standard_name = "time" ;
		time_uv:units = "seconds since 1970-01-01T00:00:00Z" ;
	char trajectory(traj_strlen) ;
		trajectory:cf_role = "trajectory_id" ;
		trajectory:comment = "A trajectory is a single deployment of a glider and may span multiple data files." ;
		trajectory:long_name = "Trajectory/Deployment Name" ;
	double u ;
		u:_FillValue = -999. ;
		u:comment = "The depth-averaged current is an estimate of the net current measured while the glider is underwater.  The value is calculated over the entire underwater segment, which may consist of 1 or more dives." ;
		u:long_name = "Depth-Averaged Eastward Sea Water Velocity" ;
		u:observation_type = "calculated" ;
		u:platform = "platform" ;
		u:standard_name = "eastward_sea_water_velocity" ;
		u:units = "m s-1" ;
		u:valid_max = 10. ;
		u:valid_min = -10. ;
	double v ;
		v:_FillValue = -999. ;
		v:comment = "The depth-averaged current is an estimate of the net current measured while the glider is underwater.  The value is calculated over the entire underwater segment, which may consist of 1 or more dives." ;
		v:long_name = "Depth-Averaged Northward Sea Water Velocity" ;
		v:observation_type = "calculated" ;
		v:platform = "platform" ;
		v:standard_name = "northward_sea_water_velocity" ;
		v:units = "m s-1" ;
		v:valid_max = 10. ;
		v:valid_min = -10. ;

// global attributes:
		:Conventions = "CF-1.6, Unidata Dataset Discovery v1.0" ;
		:Metadata_Conventions = "CF-1.6, Unidata Dataset Discovery v1.0" ;
		:acknowledgment = "This deployment supported by ..." ;
		:comment = " " ;
		:contributor_name = " " ;
		:contributor_role = " " ;
		:creator_email = " " ;
		:creator_name = " " ;
		:creator_url = " " ;
		:date_created = " " ;
		:date_issued = " " ;
		:date_modified = " " ;
		:format_version = "IOOS_Glider_NetCDF_v3.0-noqartod.nc" ;
		:history = " " ;
		:id = " " ;
		:institution = " " ;
		:ioos_regional_association = " " ;
		:keywords = "AUVS > Autonomous Underwater Vehicles, Oceans > Ocean Pressure > Water Pressure, Oceans > Ocean Temperature > Water Temperature, Oceans > Salinity/Density > Conductivity, Oceans > Salinity/Density > Density, Oceans > Salinity/Density > Salinity" ;
		:keywords_vocabulary = "GCMD Science Keywords" ;
		:license = "This data may be redistributed and used without restriction.  Data provided as is with no expressed or implied assurance of quality assurance or quality control" ;
		:metadata_link = " " ;
		:naming_authority = "edu.rutgers.marine" ;
		:platform_type = "Slocum Glider" ;
		:processing_level = " " ;
		:project = " " ;
		:publisher_email = " " ;
		:publisher_name = " " ;
		:publisher_url = " " ;
        :references = " " ;
		:sea_name = " " ;
		:source = "Observational data from a profiling glider" ;
		:standard_name_vocabulary = "CF-v25" ;
		:summary = "The Rutgers University Coastal Ocean Observation Lab has deployed autonomous underwater gliders around the world since 1990.  Gliders are small, free-swimming, unmanned vehicles that use changes in buoyancy to move vertically and horizontally through the water column in a saw-tooth pattern. They are deployed for days to several months and gather detailed information about the physical, chemical and biological processes of the world\'s The Slocum glider was designed and oceans. built by Teledyne Webb Research Corporation, Falmouth, MA, USA.  This dataset contains observational sub-surface profile data of the water-column." ;
		:title = " " ;
		:wmo_id = " " ;
}
