	double oxygen_concentration(time) ;
		oxygen_concentration:_FillValue = -999. ;
		oxygen_concentration:accuracy = " " ;
		oxygen_concentration:ancillary_variables = "oxygen_concentration_qc" ;
		oxygen_concentration:instrument = " " ;
		oxygen_concentration:long_name = "Dissolved Oxygen Concentration" ;
		oxygen_concentration:observation_type = "measured" ;
		oxygen_concentration:platform = "platform" ;
		oxygen_concentration:precision = " " ;
		oxygen_concentration:resolution = " " ;
		oxygen_concentration:standard_name = "mole_concentration_of_dissolved_molecular_oxygen_in_seawater" ;
		oxygen_concentration:units = "micromoles/L" ;
		oxygen_concentration:valid_max = 400. ;
		oxygen_concentration:valid_min = 0. ;
	byte oxygen_concentration_qc(time) ;
		oxygen_concentration_qc:_FillValue = -127b ;
		oxygen_concentration_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed not_used not_used interpolated_value missing_value" ;
		oxygen_concentration_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		oxygen_concentration_qc:long_name = "oxygen_concentration Quality Flag" ;
		oxygen_concentration_qc:standard_name = "oxygen_concentration status_flag" ;
		oxygen_concentration_qc:valid_max = 9b ;
		oxygen_concentration_qc:valid_min = 0b ;
	double oxygen_saturation(time) ;
		oxygen_saturation:_FillValue = -999. ;
		oxygen_saturation:accuracy = " " ;
		oxygen_saturation:ancillary_variables = "oxygen_saturation_qc" ;
		oxygen_saturation:instrument = " " ;
		oxygen_saturation:long_name = "Oxygen Saturation" ;
		oxygen_saturation:observation_type = "measured" ;
		oxygen_saturation:platform = "platform" ;
		oxygen_saturation:precision = " " ;
		oxygen_saturation:resolution = " " ;
		oxygen_saturation:standard_name = "fractional_saturation_of_oxygen_in_seawater" ;
		oxygen_saturation:units = "%" ;
		oxygen_saturation:valid_max = 120. ;
		oxygen_saturation:valid_min = 0. ;
	byte oxygen_saturation_qc(time) ;
		oxygen_saturation_qc:_FillValue = -127b ;
		oxygen_saturation_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed not_used not_used interpolated_value missing_value" ;
		oxygen_saturation_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		oxygen_saturation_qc:long_name = "oxygen_saturation Quality Flag" ;
		oxygen_saturation_qc:standard_name = "oxygen_saturation status_flag" ;
		oxygen_saturation_qc:valid_max = 9b ;
		oxygen_saturation_qc:valid_min = 0b ;
