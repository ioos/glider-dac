	double chlorophyll_a(time) ;
		chlorophyll_a:_FillValue = -999. ;
		chlorophyll_a:accuracy = " " ;
		chlorophyll_a:ancillary_variables = "chlorophyll_a_qc" ;
		chlorophyll_a:instrument = " " ;
		chlorophyll_a:long_name = "Chlorophyll a" ;
		chlorophyll_a:observation_type = "measured" ;
		chlorophyll_a:platform = "platform" ;
		chlorophyll_a:precision = " " ;
		chlorophyll_a:resolution = " " ;
		chlorophyll_a:standard_name = "mass_concentration_of_chlorophyll_a_in_seawater" ;
		chlorophyll_a:units = "micrograms/L" ;
		chlorophyll_a:valid_max = 40. ;
		chlorophyll_a:valid_min = 0. ;
	byte chlorophyll_a_qc(time) ;
		chlorophyll_a_qc:_FillValue = -127b ;
		chlorophyll_a_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed not_used not_used interpolated_value missing_value" ;
		chlorophyll_a_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		chlorophyll_a_qc:long_name = "chlorophyll_a Quality Flag" ;
		chlorophyll_a_qc:standard_name = "chlorophyll_a status_flag" ;
		chlorophyll_a_qc:valid_max = 9b ;
		chlorophyll_a_qc:valid_min = 0b ;
