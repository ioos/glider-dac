	double cdom(time) ;
		cdom:_FillValue = -999. ;
		cdom:accuracy = " " ;
		cdom:ancillary_variables = "cdom_qc" ;
		cdom:instrument = " " ;
		cdom:long_name = "Chromophoric Dissolved Organic Matter" ;
		cdom:observation_type = "measured" ;
		cdom:platform = "platform" ;
		cdom:precision = " " ;
		cdom:resolution = " " ;
		cdom:standard_name = " " ;
		cdom:units = "ppb" ;
		cdom:valid_max = 40. ;
		cdom:valid_min = 0. ;
	byte cdom_qc(time) ;
		cdom_qc:_FillValue = -127b ;
		cdom_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed not_used not_used interpolated_value missing_value" ;
		cdom_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		cdom_qc:long_name = "cdom Quality Flag" ;
		cdom_qc:standard_name = "cdom status_flag" ;
		cdom_qc:valid_max = 9b ;
		cdom_qc:valid_min = 0b ;
